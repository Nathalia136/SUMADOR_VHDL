library verilog;
use verilog.vl_types.all;
entity rca_4bit_vlg_vec_tst is
end rca_4bit_vlg_vec_tst;
