library verilog;
use verilog.vl_types.all;
entity DECOD7_vlg_vec_tst is
end DECOD7_vlg_vec_tst;
