library verilog;
use verilog.vl_types.all;
entity test_sum_4bits_vlg_vec_tst is
end test_sum_4bits_vlg_vec_tst;
