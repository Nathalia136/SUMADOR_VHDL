library verilog;
use verilog.vl_types.all;
entity Des_vlg_vec_tst is
end Des_vlg_vec_tst;
